module hexdecoder(c, display);
	input [4:0] c;				//4 inputs
	output [7:0] display;	//7 outputs
	
	assign display[0] = !(!c[2]&!c[0] | c[1]&!c[3] | c[1]&c[2] | c[3]&!c[0] | !c[1]&c[3]&!c[2] | !c[3]&c[2]&c[0]);
	assign display[1] = !(!c[3]&!c[2] | !c[0]&!c[2] | c[1]&c[0]&!c[3] | !c[1]&!c[0]&!c[3] | !c[1]&c[0]&c[3]);
	assign display[2] = !(c[3]&!c[2] | !c[1]&!c[3] | !c[3]&c[0] | c[2]&!c[3] | !c[1]&c[0]);
	assign display[3] = !(!c[1]&c[3] | c[1]&!c[2]&c[0] | !c[1]&c[0]&c[2] | c[2]&c[1]&!c[0] | !c[0]&!c[2]&!c[3]);
	assign display[4] = !(c[3]&c[2] | c[1]&!c[0] | c[3]&c[1] | !c[0]&!c[2]);
	assign display[5] = !(c[3]&!c[2] | !c[1]&!c[0] | c[2]&!c[0] | c[1]&c[3] | !c[3]&c[2]&!c[1]);
	assign display[6] = !(c[3]&!c[2] | c[1]&!c[0] | c[3]&c[0] | !c[3]&c[2]&!c[1] | !c[2]&c[1]);
endmodule